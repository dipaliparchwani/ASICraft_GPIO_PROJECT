`include "uvm_macros.svh"
import uvm_pkg::*;
`include "defines.sv"
`include "../sv/env/gpio_interface.sv"
`include "../sv/env/gpio_reg_interface.sv"
`include "gpio_assertion.sv"
`include "gpio_coverage.sv"
