package env_pkg; 
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import ral_pkg::*;
  import seq_pkg::*;
  `include "gpio_reg_seqr.sv"
  `include "gpio_reg_driver.sv"
  `include "gpio_reg_monitor.sv"
  `include "gpio_reg_agent.sv"
  `include "gpio_seqr.sv"
  `include "gpio_driver.sv"
  `include "gpio_monitor.sv"
  `include "gpio_agent.sv"
  `include "gpio_scoreboard.sv"
  `include "gpio_env.sv"
endpackage

