/******************************************************************************************/
/*-------------------------------------------------------------------------*/
/*PROJECT_NAME : GPIO VIP                                                  */           
/*FILE_NAME    : gpio_data_in.sv                                           */         
/*DESCRIPTION  : Read-only, Reflects the current state of the physical pins*/       
/*CREATED_ON   : 21/07/2025                                                */                                                       
/*DEVELOPER    : Dipali                                                    */
/*------------------------------------------------------------------------ */
/******************************************************************************************/
class gpio_data_in_reg extends uvm_reg;
  `uvm_object_utils(gpio_data_in_reg)

  uvm_reg_field DATA_IN;

  function new(string name = "gpio_data_in_reg");
    super.new(name,`DATA_WIDTH,UVM_NO_COVERAGE);
  endfunction

  function void build;
     DATA_IN = uvm_reg_field::type_id::create("DATA_IN");

     DATA_IN.configure( .parent(this),
                        .size(`DATA_WIDTH),
			.lsb_pos(0),
			.access("RO"),
			.volatile(1),
			.reset(0),
			.has_reset(1),
			.is_rand(0),
			.individually_accessible(1));
  endfunction
endclass
