`include "uvm_macros.svh"
import uvm_pkg::*;
`include "defines.sv"
`include "../sv/env/gpio_interface.sv"
`include "../sv/env/gpio_reg_interface.sv"
`include "gpio_assertion.sv"
package gpio_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "clk_checker.sv"
  `include "../ral/gpio_data_in_reg.sv"
  `include "../ral/gpio_data_out_reg.sv"
  `include "../ral/gpio_oe_reg.sv"
  `include "../ral/gpio_intr_mask_reg.sv"
  `include "../ral/gpio_intr_status_reg.sv"
  `include "../ral/gpio_intr_type_reg.sv"
  `include "../ral/gpio_intr_polarity_reg.sv"
  `include "../ral/gpio_dir_reg.sv"
  `include "../ral/gpio_reg_block.sv"
  `include "../seqlib/gpio_reg_transaction.sv"
  `include "../ral/gpio_adapter.sv"
  `include "../seqlib/gpio_transaction.sv"
  `include "../seqlib/reset_seq.sv"
  `include "../seqlib/in_seq.sv"
  `include "../seqlib/gpio_in_toggle_base_seq.sv"
  `include "../seqlib/gpio_in_random_seq.sv"
  `include "../seqlib/in_out_reg_seq.sv"
  `include "../seqlib/gpio_reg_reset_check_seq.sv"
  `include "../seqlib/gpio_error_seq.sv"
  `include "../seqlib/gpio_in_read_repeat_seq.sv"
  `include "../seqlib/gpio_out_write_repeat_seq.sv"
  `include "../seqlib/gpio_base_seq.sv"
  `include "../seqlib/gpio_intr_config_base_seq.sv"
  `include "../seqlib/gpio_intr_with_high_mask_seq.sv"
  `include "../seqlib/gpio_intr_with_random_mask_seq.sv"
  `include "../seqlib/gpio_intr_status_clear_seq.sv"
  `include "gpio_reg_seqr.sv"
  `include "gpio_reg_driver.sv"
  `include "gpio_reg_monitor.sv"
  `include "gpio_reg_agent.sv"
  `include "gpio_seqr.sv"
  `include "gpio_driver.sv"
  `include "gpio_monitor.sv"
  `include "gpio_agent.sv"
  `include "gpio_scoreboard.sv"
  `include "gpio_env.sv"
  `include "../../test/gpio_test.sv"
  `include "../../test/gpio_in_out_functionality_test.sv"
  `include "../../test/gpio_active_low_reset_test.sv"
  `include "../../test/gpio_error_test.sv"
  `include "../../test/gpio_in_pattern_test.sv"
  `include "../../test/gpio_in_random_test.sv"
  `include "../../test/gpio_out_random_test.sv"
  `include "../../test/gpio_intr_sanity_test.sv"
  `include "../../test/gpio_intr_random_test.sv"
  `include "../../test/gpio_intr_clear_test.sv"
endpackage
